package sreg_map_Consts;
  localparam SREG_SIZE = 4;
  localparam ADDR_SREG_AREG = 'h0;
endpackage

package enums1_Consts;
  localparam ENUMS1_SIZE = 4;
  localparam ADDR_ENUMS1_R1 = 'h0;
  localparam C_enum1_hello = 8'h0;
  localparam C_enum1_World = 8'h1;
  localparam C_enum2_hello = 1'h0;
  localparam C_enum2_world = 1'h1;
endpackage

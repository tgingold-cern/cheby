package semver1_Consts;
  localparam SEMVER1_SIZE = 4;
  localparam SEMVER1_MEMMAP_VERSION = 'h10000;
  localparam SEMVER1_IDENT = 'h12345678;
  localparam ADDR_SEMVER1_R1 = 'h0;
endpackage

package demo_all_Consts;
  localparam DEMO_ALL_SIZE = 8448;
  localparam ADDR_DEMO_ALL_REG0 = 'h0;
  localparam DEMO_ALL_REG0_FIELD00_OFFSET = 1;
  localparam DEMO_ALL_REG0_FIELD00 = 32'h2;
  localparam DEMO_ALL_REG0_FIELD01_OFFSET = 4;
  localparam DEMO_ALL_REG0_FIELD01 = 32'hf0;
  localparam DEMO_ALL_REG0_FIELD02_OFFSET = 8;
  localparam DEMO_ALL_REG0_FIELD02 = 32'h700;
  localparam ADDR_DEMO_ALL_REG1 = 'h4;
  localparam DEMO_ALL_REG1_PRESET = 32'h123;
  localparam ADDR_DEMO_ALL_REG2 = 'h8;
  localparam DEMO_ALL_REG2_FIELD10_OFFSET = 0;
  localparam DEMO_ALL_REG2_FIELD10 = 64'hffff;
  localparam DEMO_ALL_REG2_FIELD11_OFFSET = 16;
  localparam DEMO_ALL_REG2_FIELD11 = 64'hffffffffff0000;
  localparam ADDR_DEMO_ALL_BLOCK1 = 'h10;
  localparam DEMO_ALL_BLOCK1_SIZE = 16;
  localparam ADDR_DEMO_ALL_BLOCK1_B1REG0 = 'h10;
  localparam ADDR_DEMO_ALL_BLOCK1_B1REG1 = 'h14;
  localparam DEMO_ALL_BLOCK1_B1REG1_F0_OFFSET = 0;
  localparam DEMO_ALL_BLOCK1_B1REG1_F0 = 32'h1;
  localparam DEMO_ALL_BLOCK1_B1REG1_F1_OFFSET = 1;
  localparam DEMO_ALL_BLOCK1_B1REG1_F1 = 32'hfffffffe;
  localparam ADDR_DEMO_ALL_BLOCK1_B1REG2 = 'h18;
  localparam ADDR_DEMO_ALL_SUB1 = 'h20;
  localparam ADDR_MASK_DEMO_ALL_SUB1 = 'h3ff0;
  localparam DEMO_ALL_SUB1_SIZE = 16;
  localparam ADDR_DEMO_ALL_SUB2 = 'h30;
  localparam ADDR_MASK_DEMO_ALL_SUB2 = 'h3ff0;
  localparam DEMO_ALL_SUB2_SIZE = 16;
  localparam ADDR_DEMO_ALL_SUB3 = 'h1000;
  localparam ADDR_MASK_DEMO_ALL_SUB3 = 'h3000;
  localparam DEMO_ALL_SUB3_SIZE = 4096;
  localparam ADDR_DEMO_ALL_ARR1 = 'h2000;
  localparam DEMO_ALL_ARR1_SIZE = 8;
  localparam ADDR_DEMO_ALL_ARR1_0 = 'h2000;
  localparam DEMO_ALL_ARR1_0_SIZE = 4;
  localparam ADDR_DEMO_ALL_ARR1_0_AREG1 = 'h2000;
  localparam ADDR_DEMO_ALL_ARR1_1 = 'h2004;
  localparam DEMO_ALL_ARR1_1_SIZE = 4;
  localparam ADDR_DEMO_ALL_ARR1_1_AREG1 = 'h2004;
  localparam ADDR_DEMO_ALL_RAM_RO1 = 'h2080;
  localparam DEMO_ALL_RAM_RO1_SIZE = 4;
  localparam ADDR_DEMO_ALL_RAM_RO1_VALUE = 'h0;
endpackage

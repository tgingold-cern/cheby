package blkpfx_Consts is
  constant BLKPFX_SIZE : Natural := 4;
  constant ADDR_BLKPFX_REG1 : Natural := 16#0#;
end package blkpfx_Consts;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package MemMap_cregs_d8 is

  -- Ident Code
  constant C_cregs_d8_IdentCode : std_logic_vector(7 downto 0) := X"FF";

  -- Memory Map Version
  constant C_cregs_d8_MemMapVersion : std_logic_vector(31 downto 0) := X"0133A207";--20161031
  -- Register Addresses : Memory Map
  constant C_Reg_cregs_d8_test1_3 : std_logic_vector(19 downto 0) := "00000000000000000000";-- : Word address : "0" & X"00000"; Byte Address : X"00000"
  constant C_Reg_cregs_d8_test1_2 : std_logic_vector(19 downto 0) := "00000000000000000001";-- : Word address : "0" & X"00001"; Byte Address : X"00002"
  constant C_Reg_cregs_d8_test1_1 : std_logic_vector(19 downto 0) := "00000000000000000010";-- : Word address : "0" & X"00002"; Byte Address : X"00004"
  constant C_Reg_cregs_d8_test1_0 : std_logic_vector(19 downto 0) := "00000000000000000011";-- : Word address : "0" & X"00003"; Byte Address : X"00006"
  constant C_Reg_cregs_d8_test2_3 : std_logic_vector(19 downto 0) := "00000000000000000100";-- : Word address : "0" & X"00004"; Byte Address : X"00008"
  constant C_Reg_cregs_d8_test2_2 : std_logic_vector(19 downto 0) := "00000000000000000101";-- : Word address : "0" & X"00005"; Byte Address : X"0000a"
  constant C_Reg_cregs_d8_test2_1 : std_logic_vector(19 downto 0) := "00000000000000000110";-- : Word address : "0" & X"00006"; Byte Address : X"0000c"
  constant C_Reg_cregs_d8_test2_0 : std_logic_vector(19 downto 0) := "00000000000000000111";-- : Word address : "0" & X"00007"; Byte Address : X"0000e"
  constant C_Reg_cregs_d8_test3_3 : std_logic_vector(19 downto 0) := "00000000000000001000";-- : Word address : "0" & X"00008"; Byte Address : X"00010"
  constant C_Reg_cregs_d8_test3_2 : std_logic_vector(19 downto 0) := "00000000000000001001";-- : Word address : "0" & X"00009"; Byte Address : X"00012"
  constant C_Reg_cregs_d8_test3_1 : std_logic_vector(19 downto 0) := "00000000000000001010";-- : Word address : "0" & X"0000a"; Byte Address : X"00014"
  constant C_Reg_cregs_d8_test3_0 : std_logic_vector(19 downto 0) := "00000000000000001011";-- : Word address : "0" & X"0000b"; Byte Address : X"00016"
  constant C_Reg_cregs_d8_test4_3 : std_logic_vector(19 downto 0) := "00000000000000001100";-- : Word address : "0" & X"0000c"; Byte Address : X"00018"
  constant C_Reg_cregs_d8_test4_2 : std_logic_vector(19 downto 0) := "00000000000000001101";-- : Word address : "0" & X"0000d"; Byte Address : X"0001a"
  constant C_Reg_cregs_d8_test4_1 : std_logic_vector(19 downto 0) := "00000000000000001110";-- : Word address : "0" & X"0000e"; Byte Address : X"0001c"
  constant C_Reg_cregs_d8_test4_0 : std_logic_vector(19 downto 0) := "00000000000000001111";-- : Word address : "0" & X"0000f"; Byte Address : X"0001e"
  constant C_Reg_cregs_d8_test5_3 : std_logic_vector(19 downto 0) := "00000000000000010000";-- : Word address : "0" & X"00010"; Byte Address : X"00020"
  constant C_Reg_cregs_d8_test5_2 : std_logic_vector(19 downto 0) := "00000000000000010001";-- : Word address : "0" & X"00011"; Byte Address : X"00022"
  constant C_Reg_cregs_d8_test5_1 : std_logic_vector(19 downto 0) := "00000000000000010010";-- : Word address : "0" & X"00012"; Byte Address : X"00024"
  constant C_Reg_cregs_d8_test5_0 : std_logic_vector(19 downto 0) := "00000000000000010011";-- : Word address : "0" & X"00013"; Byte Address : X"00026"
  constant C_Reg_cregs_d8_test6_3 : std_logic_vector(19 downto 0) := "00000000000000010100";-- : Word address : "0" & X"00014"; Byte Address : X"00028"
  constant C_Reg_cregs_d8_test6_2 : std_logic_vector(19 downto 0) := "00000000000000010101";-- : Word address : "0" & X"00015"; Byte Address : X"0002a"
  constant C_Reg_cregs_d8_test6_1 : std_logic_vector(19 downto 0) := "00000000000000010110";-- : Word address : "0" & X"00016"; Byte Address : X"0002c"
  constant C_Reg_cregs_d8_test6_0 : std_logic_vector(19 downto 0) := "00000000000000010111";-- : Word address : "0" & X"00017"; Byte Address : X"0002e"
  constant C_Reg_cregs_d8_test7_3 : std_logic_vector(19 downto 0) := "00000000000000011000";-- : Word address : "0" & X"00018"; Byte Address : X"00030"
  constant C_Reg_cregs_d8_test7_2 : std_logic_vector(19 downto 0) := "00000000000000011001";-- : Word address : "0" & X"00019"; Byte Address : X"00032"
  constant C_Reg_cregs_d8_test7_1 : std_logic_vector(19 downto 0) := "00000000000000011010";-- : Word address : "0" & X"0001a"; Byte Address : X"00034"
  constant C_Reg_cregs_d8_test7_0 : std_logic_vector(19 downto 0) := "00000000000000011011";-- : Word address : "0" & X"0001b"; Byte Address : X"00036"
  constant C_Reg_cregs_d8_test8_3 : std_logic_vector(19 downto 0) := "00000000000000011100";-- : Word address : "0" & X"0001c"; Byte Address : X"00038"
  constant C_Reg_cregs_d8_test8_2 : std_logic_vector(19 downto 0) := "00000000000000011101";-- : Word address : "0" & X"0001d"; Byte Address : X"0003a"
  constant C_Reg_cregs_d8_test8_1 : std_logic_vector(19 downto 0) := "00000000000000011110";-- : Word address : "0" & X"0001e"; Byte Address : X"0003c"
  constant C_Reg_cregs_d8_test8_0 : std_logic_vector(19 downto 0) := "00000000000000011111";-- : Word address : "0" & X"0001f"; Byte Address : X"0003e"

  -- Register Auto Clear Masks : Memory Map
  constant C_ACM_cregs_d8_test1_3 : std_logic_vector(15 downto 12) := "0000";-- : Value : X"0"
  constant C_ACM_cregs_d8_test1_2 : std_logic_vector(11 downto 8) := "0000";-- : Value : X"0"
  constant C_ACM_cregs_d8_test1_1 : std_logic_vector(7 downto 4) := "0000";-- : Value : X"0"
  constant C_ACM_cregs_d8_test1_0 : std_logic_vector(3 downto 0) := "0000";-- : Value : X"0"
  constant C_ACM_cregs_d8_test2_3 : std_logic_vector(15 downto 12) := "0000";-- : Value : X"0"
  constant C_ACM_cregs_d8_test2_2 : std_logic_vector(11 downto 8) := "0000";-- : Value : X"0"
  constant C_ACM_cregs_d8_test2_1 : std_logic_vector(7 downto 4) := "0000";-- : Value : X"0"
  constant C_ACM_cregs_d8_test2_0 : std_logic_vector(3 downto 0) := "0000";-- : Value : X"0"
  constant C_ACM_cregs_d8_test3_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test3_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test3_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test3_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test4_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test4_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test4_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test4_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test5_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test5_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test5_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test5_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test6_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test6_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test6_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test6_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test7_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test7_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test7_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test7_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test8_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test8_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test8_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_ACM_cregs_d8_test8_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"

  -- Register Preset Masks : Memory Map
  constant C_PSM_cregs_d8_test1_3 : std_logic_vector(15 downto 12) := "0000";-- : Value : X"0"
  constant C_PSM_cregs_d8_test1_2 : std_logic_vector(11 downto 8) := "0000";-- : Value : X"0"
  constant C_PSM_cregs_d8_test1_1 : std_logic_vector(7 downto 4) := "0000";-- : Value : X"0"
  constant C_PSM_cregs_d8_test1_0 : std_logic_vector(3 downto 0) := "0000";-- : Value : X"0"
  constant C_PSM_cregs_d8_test2_3 : std_logic_vector(15 downto 12) := "0000";-- : Value : X"0"
  constant C_PSM_cregs_d8_test2_2 : std_logic_vector(11 downto 8) := "0000";-- : Value : X"0"
  constant C_PSM_cregs_d8_test2_1 : std_logic_vector(7 downto 4) := "0000";-- : Value : X"0"
  constant C_PSM_cregs_d8_test2_0 : std_logic_vector(3 downto 0) := "0000";-- : Value : X"0"
  constant C_PSM_cregs_d8_test3_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test3_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test3_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test3_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test4_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test4_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test4_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test4_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test5_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test5_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test5_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test5_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test6_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test6_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test6_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test6_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test7_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test7_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test7_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test7_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test8_3 : std_logic_vector(31 downto 24) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test8_2 : std_logic_vector(23 downto 16) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test8_1 : std_logic_vector(15 downto 8) := "00000000";-- : Value : X"00"
  constant C_PSM_cregs_d8_test8_0 : std_logic_vector(7 downto 0) := "00000000";-- : Value : X"00"

  -- CODE FIELDS
  -- Memory Data : Memory Map
  -- Submap Addresses : Memory Map
end MemMap_cregs_d8;

library ieee;
use ieee.std_logic_1164.all;

package top_Consts is
  constant TOP_SIZE : Natural := 32;
  constant ADDR_TOP_ARRAY_OF_SUBMAPS : Natural := 16#0#;
  constant TOP_ARRAY_OF_SUBMAPS_SIZE : Natural := 32;
  constant ADDR_TOP_ARRAY_OF_SUBMAPS_0 : Natural := 16#0#;
  constant TOP_ARRAY_OF_SUBMAPS_0_SIZE : Natural := 4;
  constant ADDR_TOP_ARRAY_OF_SUBMAPS_0_SUBMAP : Natural := 16#0#;
  constant ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_0_SUBMAP : Natural := 16#1c#;
  constant TOP_ARRAY_OF_SUBMAPS_0_SUBMAP_SIZE : Natural := 4;
  constant ADDR_TOP_ARRAY_OF_SUBMAPS_1 : Natural := 16#4#;
  constant TOP_ARRAY_OF_SUBMAPS_1_SIZE : Natural := 4;
  constant ADDR_TOP_ARRAY_OF_SUBMAPS_1_SUBMAP : Natural := 16#4#;
  constant ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_1_SUBMAP : Natural := 16#1c#;
  constant TOP_ARRAY_OF_SUBMAPS_1_SUBMAP_SIZE : Natural := 4;
  constant ADDR_TOP_ARRAY_OF_SUBMAPS_2 : Natural := 16#8#;
  constant TOP_ARRAY_OF_SUBMAPS_2_SIZE : Natural := 4;
  constant ADDR_TOP_ARRAY_OF_SUBMAPS_2_SUBMAP : Natural := 16#8#;
  constant ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_2_SUBMAP : Natural := 16#1c#;
  constant TOP_ARRAY_OF_SUBMAPS_2_SUBMAP_SIZE : Natural := 4;
  constant ADDR_TOP_ARRAY_OF_SUBMAPS_3 : Natural := 16#c#;
  constant TOP_ARRAY_OF_SUBMAPS_3_SIZE : Natural := 4;
  constant ADDR_TOP_ARRAY_OF_SUBMAPS_3_SUBMAP : Natural := 16#c#;
  constant ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_3_SUBMAP : Natural := 16#1c#;
  constant TOP_ARRAY_OF_SUBMAPS_3_SUBMAP_SIZE : Natural := 4;
  constant ADDR_TOP_ARRAY_OF_SUBMAPS_4 : Natural := 16#10#;
  constant TOP_ARRAY_OF_SUBMAPS_4_SIZE : Natural := 4;
  constant ADDR_TOP_ARRAY_OF_SUBMAPS_4_SUBMAP : Natural := 16#10#;
  constant ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_4_SUBMAP : Natural := 16#1c#;
  constant TOP_ARRAY_OF_SUBMAPS_4_SUBMAP_SIZE : Natural := 4;
end package top_Consts;

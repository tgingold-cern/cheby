library ieee;
use ieee.std_logic_1164.all;

package sreg_map_Consts is
  constant SREG_SIZE : Natural := 4;
  constant ADDR_SREG_AREG : Natural := 16#0#;
end package sreg_map_Consts;

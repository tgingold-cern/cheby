package pkg_top_consts;
  localparam TOP_SIZE = 32;
  localparam ADDR_TOP_ARRAY_OF_SUBMAPS = 'h0;
  localparam ADDR_MASK_TOP_ARRAY_OF_SUBMAPS = 'h0;
  localparam ADDR_FMASK_TOP_ARRAY_OF_SUBMAPS = 'h0;
  localparam TOP_ARRAY_OF_SUBMAPS_SIZE = 32;
  localparam ADDR_TOP_ARRAY_OF_SUBMAPS_0 = 'h0;
  localparam ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_0 = 'h1c;
  localparam ADDR_FMASK_TOP_ARRAY_OF_SUBMAPS_0 = 'h1c;
  localparam TOP_ARRAY_OF_SUBMAPS_0_SIZE = 4;
  localparam ADDR_TOP_ARRAY_OF_SUBMAPS_0_SUBMAP = 'h0;
  localparam ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_0_SUBMAP = 'h1c;
  localparam ADDR_FMASK_TOP_ARRAY_OF_SUBMAPS_0_SUBMAP = 'h1c;
  localparam TOP_ARRAY_OF_SUBMAPS_0_SUBMAP_SIZE = 4;
  localparam ADDR_TOP_ARRAY_OF_SUBMAPS_1 = 'h4;
  localparam ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_1 = 'h1c;
  localparam ADDR_FMASK_TOP_ARRAY_OF_SUBMAPS_1 = 'h1c;
  localparam TOP_ARRAY_OF_SUBMAPS_1_SIZE = 4;
  localparam ADDR_TOP_ARRAY_OF_SUBMAPS_1_SUBMAP = 'h4;
  localparam ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_1_SUBMAP = 'h1c;
  localparam ADDR_FMASK_TOP_ARRAY_OF_SUBMAPS_1_SUBMAP = 'h1c;
  localparam TOP_ARRAY_OF_SUBMAPS_1_SUBMAP_SIZE = 4;
  localparam ADDR_TOP_ARRAY_OF_SUBMAPS_2 = 'h8;
  localparam ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_2 = 'h1c;
  localparam ADDR_FMASK_TOP_ARRAY_OF_SUBMAPS_2 = 'h1c;
  localparam TOP_ARRAY_OF_SUBMAPS_2_SIZE = 4;
  localparam ADDR_TOP_ARRAY_OF_SUBMAPS_2_SUBMAP = 'h8;
  localparam ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_2_SUBMAP = 'h1c;
  localparam ADDR_FMASK_TOP_ARRAY_OF_SUBMAPS_2_SUBMAP = 'h1c;
  localparam TOP_ARRAY_OF_SUBMAPS_2_SUBMAP_SIZE = 4;
  localparam ADDR_TOP_ARRAY_OF_SUBMAPS_3 = 'hc;
  localparam ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_3 = 'h1c;
  localparam ADDR_FMASK_TOP_ARRAY_OF_SUBMAPS_3 = 'h1c;
  localparam TOP_ARRAY_OF_SUBMAPS_3_SIZE = 4;
  localparam ADDR_TOP_ARRAY_OF_SUBMAPS_3_SUBMAP = 'hc;
  localparam ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_3_SUBMAP = 'h1c;
  localparam ADDR_FMASK_TOP_ARRAY_OF_SUBMAPS_3_SUBMAP = 'h1c;
  localparam TOP_ARRAY_OF_SUBMAPS_3_SUBMAP_SIZE = 4;
  localparam ADDR_TOP_ARRAY_OF_SUBMAPS_4 = 'h10;
  localparam ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_4 = 'h1c;
  localparam ADDR_FMASK_TOP_ARRAY_OF_SUBMAPS_4 = 'h1c;
  localparam TOP_ARRAY_OF_SUBMAPS_4_SIZE = 4;
  localparam ADDR_TOP_ARRAY_OF_SUBMAPS_4_SUBMAP = 'h10;
  localparam ADDR_MASK_TOP_ARRAY_OF_SUBMAPS_4_SUBMAP = 'h1c;
  localparam ADDR_FMASK_TOP_ARRAY_OF_SUBMAPS_4_SUBMAP = 'h1c;
  localparam TOP_ARRAY_OF_SUBMAPS_4_SUBMAP_SIZE = 4;
endpackage

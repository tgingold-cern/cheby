package fid_top_axi_Consts;
  localparam FID_TOP_AXI_MEMMAP_VERSION = 'h100;
  localparam ADDR_FID_TOP_AXI_IP = 'h0;
  localparam ADDR_MASK_FID_TOP_AXI_IP = 'h0;
  localparam ADDR_FMASK_FID_TOP_AXI_IP = 'h0;
  localparam FID_TOP_AXI_IP_SIZE = 4;
endpackage

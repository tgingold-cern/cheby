package semver1_Consts is
  constant SEMVER1_SIZE : Natural := 4;
  constant SEMVER1_VERSION : Natural := 16#10000#;
  constant ADDR_SEMVER1_R1 : Natural := 16#0#;
end package semver1_Consts;

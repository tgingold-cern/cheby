package memwide_ua_Consts;
  localparam MEMWIDE_UA_SIZE = 256;
  localparam ADDR_MEMWIDE_UA_REGA = 'h0;
  localparam ADDR_MEMWIDE_UA_REGA_FIELD0 = 'h0;
  localparam MEMWIDE_UA_REGA_FIELD0_OFFSET = 1;
  localparam MEMWIDE_UA_REGA_FIELD0 = 32'h2;
  localparam ADDR_MEMWIDE_UA_TS = 'h80;
  localparam MEMWIDE_UA_TS_SIZE = 16;
  localparam ADDR_MEMWIDE_UA_TS_RISE_SEC = 'h0;
  localparam ADDR_MEMWIDE_UA_TS_RISE_NS = 'h4;
  localparam ADDR_MEMWIDE_UA_TS_FALL_SEC = 'h8;
endpackage

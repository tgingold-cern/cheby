package blkpfx_Consts;
  localparam BLKPFX_SIZE = 4;
  localparam ADDR_BLKPFX_REG1 = 'h0;
endpackage

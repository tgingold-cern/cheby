package const_range_Consts;
  localparam CONST_RANGE_SIZE = 20;
  localparam ADDR_CONST_RANGE_LARGE_VAL_0 = 'h0;
  localparam CONST_RANGE_LARGE_VAL_0_PRESET = 32'hf38243bb;
  localparam ADDR_CONST_RANGE_LARGE_VAL_1 = 'h4;
  localparam CONST_RANGE_LARGE_VAL_1_PRESET = 32'hfffffff7;
  localparam ADDR_CONST_RANGE_SUPER_LARGE_VAL = 'h8;
  localparam CONST_RANGE_SUPER_LARGE_VAL_PRESET = 64'h818734fa9b1e0cf4;
  localparam ADDR_CONST_RANGE_SMALL_VAL = 'h10;
  localparam CONST_RANGE_SMALL_VAL_PRESET = 32'h1;
endpackage

package same_label_reg_Consts;
  localparam SAME_LABEL_REG_SIZE = 16;
  localparam ADDR_SAME_LABEL_REG_NO_FIELDS = 'h0;
  localparam SAME_LABEL_REG_NO_FIELDS_PRESET = 8'h20;
  localparam ADDR_SAME_LABEL_REG_SAME_NAME = 'h4;
  localparam SAME_LABEL_REG_SAME_NAME_WIDTH = 1;
  localparam SAME_LABEL_REG_SAME_NAME_OFFSET = 0;
  localparam SAME_LABEL_REG_SAME_NAME = 32'h1;
  localparam ADDR_SAME_LABEL_REG_SAME_NAME_MULTI = 'h8;
  localparam SAME_LABEL_REG_SAME_NAME_MULTI_WIDTH = 12;
  localparam SAME_LABEL_REG_SAME_NAME_MULTI_OFFSET = 0;
  localparam SAME_LABEL_REG_SAME_NAME_MULTI = 32'hfff;
  localparam ADDR_SAME_LABEL_REG_NOT_SAME_REG = 'hc;
  localparam ADDR_SAME_LABEL_REG_NOT_SAME = 'hc;
  localparam SAME_LABEL_REG_NOT_SAME_WIDTH = 1;
  localparam SAME_LABEL_REG_NOT_SAME_OFFSET = 0;
  localparam SAME_LABEL_REG_NOT_SAME = 32'h1;
endpackage

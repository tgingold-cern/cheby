package enums2_Consts;
  localparam ENUMS2_SIZE = 4;
  localparam ADDR_ENUMS2_R1 = 'h0;
  localparam ENUMS2_R1_F1_OFFSET = 0;
  localparam ENUMS2_R1_F1 = 32'hff;
  localparam C_enum1_hello = 8'h0;
  localparam C_enum1_World = 8'h1;
  localparam C_enum2_hello = 1'h0;
  localparam C_enum2_world = 1'h1;
endpackage

package semver1_Consts;
  localparam SEMVER1_SIZE = 4;
  localparam SEMVER1_VERSION = 'h10000;
  localparam ADDR_SEMVER1_R1 = 'h0;
endpackage
